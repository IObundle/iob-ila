//data and address widths
`define ILA_RDATA_W 32
`define ILA_WDATA_W 16
`define ILA_ADDR_W 3

