`ifndef DATA_W
 `define DATA_W 32
`endif

//data and address widths
`define ILA_RDATA_W 32
`define ILA_WDATA_W 32
`define ILA_ADDR_W 4

`define ILA_MAX_TRIGGERS        32
`define ILA_MAX_SAMPLES_W       16
`define ILA_MAX_SIGNAL_SELECT_W 4

`define ILA_SINGLE_TYPE     0
`define ILA_CONTINUOUS_TYPE 1

`define ILA_REDUCE_OR  0
`define ILA_REDUCE_AND 1
