`define CEIL_DIV(A, B) (A % B == 0 ? (A / B) : ((A/B) + 1))
