//data and address widths
`define ILA_RDATA_W 32
`define ILA_WDATA_W 16
`define ILA_ADDR_W 3

`define ILA_SIGNAL_W            32

`define ILA_MAX_TRIGGERS        8
`define ILA_MAX_SAMPLES_W       12
`define ILA_MAX_SIGNAL_SELECT_W 1

`define ILA_SINGLE_TYPE     1'b0
`define ILA_CONTINUOUS_TYPE 1'b1

`define ILA_REDUCE_OR  1'b0
`define ILA_REDUCE_AND 1'b1
